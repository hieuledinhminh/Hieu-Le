module alu_tb;
   reg	 [3:0] a;
   reg	 [3:0] b;
   reg	 [2:0] op;
   reg	 rst_n;
   reg	 clk;
   reg	 [3:0] result;
   reg	 carry;
   synth_wrapper alu(
	.a(a),
	.b(b),
        .rst_n(rst_n),
        .clk(clk),
	.op(op),
	.result(result),
	.carry(carry)
   );
initial begin
#0 clk=1'b0;
end
always #50 clk=~clk;

initial begin

#0
	rst_n = 1'b1; 
	a = 4'b1111;
	b = 4'b0000;
	op = 3'b111; 
#500	
	a = 4'b1010;
	b = 4'b1111;
	op = 3'b001; 
#1000	
	op = 4'b111;
	a = 4'b1111; 
	b = 4'b0010;
#1500	
	rst_n = 1'b0;
	a = 4'b1111;
	b = 4'b0000;
	op = 3'b111;
#2000	
	a = 4'b1111;
	b = 4'b0001;
	op = 3'b111;
#2500	
	a = 4'b1111;
	b = 4'b0010;
	op = 3'b111;
#3000	
	a = 4'b1111;
	b = 4'b0011;
	op = 3'b111;
#3500	
	a = 4'b1111;
	b = 4'b0100;
	op = 3'b111;
#4000	
	a = 4'b1111;
	b = 4'b0101;
	op = 3'b111;
#4500	
	a = 4'b1111;
	b = 4'b0000;
	op = 3'b110;
#5000	
	a = 4'b1111;
	b = 4'b0001;
	op = 3'b110;
#5500	
	a = 4'b1111;
	b = 4'b0010;
	op = 3'b110;
#6000	
	a = 4'b1111;
	b = 4'b0011;
	op = 3'b110;
#6500	
	a = 4'b1111;
	b = 4'b0100;
	op = 3'b110;
#7000	
	a = 4'b1111;
	b = 4'b0101;
	op = 3'b110;
#7500	
	a = 4'b1111;
	b = 4'b0101;
	op = 3'b110;
#8000	
	rst_n = 1'b1;
	a = 4'b1010;
	b = 4'b0101;
	op = 3'b110;
#8500	
	rst_n = 1'b1;
	a = 4'b0101;
	b = 4'b0101;
	op = 3'b110;
#9000	
	rst_n = 1'b1;
	a = 4'b0110;
	b = 4'b0101;
	op = 3'b110;
#9500	
	rst_n = 1'b1;
	a = 4'b1001;
	b = 4'b0101;
	op = 3'b110;
#10000	
	rst_n = 1'b1;
	a = 4'b0000;
	b = 4'b0101;
	op = 3'b110;
#10500	
	rst_n = 1'b0;
	a = 4'b0000;
	b = 4'b0101;
	op = 3'b101;
#11000	
	a = 4'b1010;
	b = 4'b0101;
	op = 3'b101;
#11500	
	a = 4'b1100;
	b = 4'b0110;
	op = 3'b101;
#12000	
	a = 4'b1100;
	b = 4'b0110;
	op = 3'b100;
#12500	
	a = 4'b0000;
	b = 4'b0110;
	op = 3'b100;
#13000	
	a = 4'b1111;
	b = 4'b0110;
	op = 3'b100;
#13500	
	a = 4'b1010;
	b = 4'b0110;
	op = 3'b100;
#14000	
	a = 4'b1100;
	b = 4'b0110;
	op = 3'b010;
#14500	
	a = 4'b0000;
	b = 4'b0110;
	op = 3'b010;
#15000	
	a = 4'b1111;
	b = 4'b0110;
	op = 3'b010;
#15500	
	a = 4'b1010;
	b = 4'b0110;
	op = 3'b001;
#16000	
	a = 4'b1010;
	b = 4'b0110;
	op = 3'b001;
#16500	
	a = 4'b0010;
	b = 4'b0110;
	op = 3'b001;
#17000	
	a = 4'b1110;
	b = 4'b0110;
	op = 3'b001;
#17500	
	a = 4'b1010;
	b = 4'b1010;
	op = 3'b001;
#18000	
	a = 4'b0000;
	b = 4'b1010;
	op = 3'b010;
#18500	
	a = 4'b0000;
	b = 4'b0101;
	op = 3'b000;
#19000	
	a = 4'b1100;
	b = 4'b0110;
	op = 3'b000;
#19500	
	a = 4'b0000;
	b = 4'b0110;
	op = 3'b000;
#20000	
	a = 4'b1111;
	b = 4'b0110;
	op = 3'b000;
#20500	
	a = 4'b1010;
	b = 4'b0110;
	op = 3'b000;
#21000	
	a = 4'b1010;
	b = 4'b0110;
	op = 3'b000;
#21500	
	a = 4'b0010;
	b = 4'b0110;
	op = 3'b000;
#22000	
	a = 4'b1110;
	b = 4'b0110;
	op = 3'b000;
#22500	
	a = 4'b1010;
	b = 4'b1010;
	op = 3'b000;
#23000	
	a = 4'b0000;
	b = 4'b1010;
	op = 3'b000;
#23500
	a = 4'b1010;
	b = 4'b0101;
	op = 3'b011;
#24000
	a = 4'b0110;
	b = 4'b1100;
	op = 3'b011;
#24500	
	a = 4'b1110;
	b = 4'b1100;
	op = 3'b011;
#25000	
	a = 4'b0001;
	b = 4'b1111;
	op = 3'b011;
end
endmodule 
